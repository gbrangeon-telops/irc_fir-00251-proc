-------------------------------------------------------------------------------
--
-- Title       : Stim
-- Design      : Line_Buffer
-- Author      : ETD
-- Company     : Telops
--
-------------------------------------------------------------------------------
--
-- File        : D:\Telops\2020-08-08 Line Buffer\Simulation\Line_buffer\src\Stim.vhd
-- Generated   : Mon Aug 31 14:28:25 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : Fichier de stimulation et de vérification pour le testbench du line buffer
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use ieee.numeric_std.all;
use work.tel2000.all;	
library std;
use std.textio.all;
use ieee.std_logic_textio.all;



entity scd_proxy2_dsync_tb is
	--port();
end scd_proxy2_dsync_tb;


architecture scd_proxy2_dsync_tb of scd_proxy2_dsync_tb is	

function hex_string_to_std_logic_vector(s: string)	return std_logic_vector is
	variable slv : std_logic_vector((s'high-s'low+1)*4-1 downto 0);
	variable k : integer;
begin
	k := s'high-s'low;
	for i in s'range loop
		case s(i) is
			when '0' =>
				slv(k*4+3 downto k*4) := x"0";
			when '1' =>
				slv(k*4+3 downto k*4) := x"1";
			when '2' =>
				slv(k*4+3 downto k*4) := x"2";
			when '3' =>
				slv(k*4+3 downto k*4) := x"3";
			when '4' =>
				slv(k*4+3 downto k*4) := x"4";
			when '5' =>
				slv(k*4+3 downto k*4) := x"5";
			when '6' =>
				slv(k*4+3 downto k*4) := x"6";
			when '7' =>
				slv(k*4+3 downto k*4) := x"7";
			when '8' =>
				slv(k*4+3 downto k*4) := x"8";
			when '9' =>
				slv(k*4+3 downto k*4) := x"9";
			when 'A' =>
				slv(k*4+3 downto k*4) := x"A";
			when 'B' =>
				slv(k*4+3 downto k*4) := x"B";
			when 'C' =>
				slv(k*4+3 downto k*4) := x"C";
			when 'D' =>
				slv(k*4+3 downto k*4) := x"D";
			when 'E' =>
				slv(k*4+3 downto k*4) := x"E";
			when 'F' =>
				slv(k*4+3 downto k*4) := x"F";
			when 'U' =>
				slv(k*4+3 downto k*4) := "UUUU";
			when 'X' =>
				slv(k*4+3 downto k*4) := "XXXX"; 
			when 'Z' =>
				slv(k*4+3 downto k*4) := "ZZZZ";
			when 'W' =>
				slv(k*4+3 downto k*4) := "WWWW";
			when 'L' =>
				slv(k*4+3 downto k*4) := "LLLL";
			when 'H' =>
				slv(k*4+3 downto k*4) := "HHHH"; 
			when '-' =>
				slv(k*4+3 downto k*4) := "----"; 
			when others =>
				slv(k*4+3 downto k*4) := "XXXX";
		end case;	
		k := k-1;
	end loop;	 
	return slv;
end hex_string_to_std_logic_vector;

component scd_proxy2_dsync
   port(
		CLK_CH0 : in std_logic;
      CLK_CH1 : in std_logic;
      D_CLK : in std_logic;
		ARESET : in std_logic;
		 
		CH0_DATA : in std_logic_vector(31 downto 0);
      CH0_DVAL : in std_logic;
      CH1_DATA : in std_logic_vector(31 downto 0);
      CH1_DVAL : in std_logic;
      
      QUAD_DATA_OUT : out std_logic_vector(71 downto 0);
	   QUAD_DVAL : out std_logic
      );
end component;

signal datatosave : std_logic_vector(63 downto 0);

file stimulus_image0 : text;
file stimulus_image1 : text;
file stimulus_start_up : text;

constant clk_period : time := 10 ns;
signal clk_i : std_logic;
signal ARESET : std_logic;
signal ch_data0 : std_logic_vector(31 downto 0);
signal ch_dval0 : std_logic;
signal ch_data1 : std_logic_vector(31 downto 0);
signal ch_dval1 : std_logic;
signal quad_data_out : std_logic_vector(71 downto 0);
signal quad_dval : std_logic;

begin

	--Clock 100Mhz definition
   clk_100Mhz_process : process
   begin 
      clk_i <= '0';
      wait for clk_period/2;
      clk_i <= '1';
      wait for clk_period/2;
   end process;
   
   --The format of stimulus_lineX needs to be 4 hex per line
	read_image_process0 : process
		variable l : line;
		variable s : string(1 to 8);
	begin
	  
      ch_dval0 <= '0';
      
      wait for clk_period * 50;
      
      --Read the image in an infinite loop like the detector would
      --Only one image is read in a loop
      while true loop
         file_open(stimulus_image0, "D:\Telops\FIR-00251-Proc\src\bb1920_serdes\SIM\Dsync0.txt",  read_mode);
         while not endfile(stimulus_image0) loop
            wait until rising_edge(clk_i);	
            readline(stimulus_image0,l);
            read(l,s);
            ch_data0 <= hex_string_to_std_logic_vector(s); 
            ch_dval0 <= '1';
         end loop;		
         file_close(stimulus_image0);
         ch_dval0 <= '0';
		end loop;
      
      wait;
	end process read_image_process0;
   
      --The format of stimulus_lineX needs to be 4 hex per line
	read_image_process1 : process
		variable l : line;
		variable s : string(1 to 8);
	begin
      
      ch_dval1 <= '0';
	  
      wait for clk_period * 50;
      
      --Read the image in an infinite loop like the detector would
      --Only one image is read in a loop
      while true loop
         file_open(stimulus_image1, "D:\Telops\FIR-00251-Proc\src\bb1920_serdes\SIM\Dsync1.txt",  read_mode);
         while not endfile(stimulus_image1) loop
            wait until rising_edge(clk_i);	
            readline(stimulus_image1,l);
            read(l,s);
            ch_data1 <= hex_string_to_std_logic_vector(s);  
            ch_dval1 <= '1';
         end loop;		
         file_close(stimulus_image1);
         ch_dval1 <= '0';
		end loop;
      
      wait;
	end process read_image_process1;
   
   gen_stim : process
   begin
      ARESET <= '1';
      
      wait for clk_period * 5;
      
      ARESET <= '0';
      
      wait;
   end process;
   
   uut: scd_proxy2_dsync
   port map(
	  CLK_CH0 => clk_i,
      CLK_CH1 => clk_i,
      D_CLK => clk_i,
	  ARESET => ARESET,
		 
      CH0_DATA => ch_data0,
      CH0_DVAL => ch_dval0,
      CH1_DATA => ch_data1,
      CH1_DVAL => ch_dval1,
      
      QUAD_DATA_OUT => quad_data_out,
	   QUAD_DVAL => quad_dval);

end scd_proxy2_dsync_tb;
