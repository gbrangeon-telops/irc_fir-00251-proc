-----------------------------------------------------------------
--!   @file mb_model_wrapper.vhd
--!   @brief Wrapper for the microblaze model.
--!   @details This component map different AXI4Lite Port.
--!
--!   $Rev$
--!   $Author$
--!   $Date$
--!   $Id$
--!   $URL$
------------------------------------------------------------------

--!   Use IEEE standard library.
library IEEE;
--!   Use logic elements package from IEEE library.
use IEEE.STD_LOGIC_1164.all; 
--!   Use TEL2000 package package from work library. 
use work.TEL2000.all;

entity mb_model_wrapper is
port(

   ACLK : in std_logic; --! Clock for core logic
   ARESETN : in std_logic; --! Reset active low for core logic
   
   GPIO_MOSI : out t_axi4_lite_mosi;
   GPIO_MISO : in t_axi4_lite_miso;

   USB_UART_MOSI : out t_axi4_lite_mosi;
   USB_UART_MISO : in t_axi4_lite_miso;

   CLINK_UART_MOSI : out t_axi4_lite_mosi;
   CLINK_UART_MISO : in t_axi4_lite_miso;
   
   FPGA_UART_MOSI : out t_axi4_lite_mosi;
   FPGA_UART_MISO : in t_axi4_lite_miso;
   
   OEM_UART_MOSI : out t_axi4_lite_mosi;
   OEM_UART_MISO : in t_axi4_lite_miso;
   
   PLEORA_UART_MOSI : out t_axi4_lite_mosi;
   PLEORA_UART_MISO : in t_axi4_lite_miso;
   
   XADC_MOSI : out t_axi4_lite_mosi;
   XADC_MISO : in t_axi4_lite_miso;

   INTC_MOSI : out t_axi4_lite_mosi;
   INTC_MISO : in t_axi4_lite_miso;

   AEC_CTRL_MOSI : out t_axi4_lite_mosi;
   AEC_CTRL_MISO : in t_axi4_lite_miso;
   
   BPR_CTRL_MOSI : out t_axi4_lite_mosi;
   BPR_CTRL_MISO : in t_axi4_lite_miso;

   CAL_CTRL_MOSI : out t_axi4_lite_mosi;
   CAL_CTRL_MISO : in t_axi4_lite_miso;
   
   EXPTIME_CTRL_MOSI : out t_axi4_lite_mosi;
   EXPTIME_CTRL_MISO : in t_axi4_lite_miso;
   
   FPA_CTRL_MOSI : out t_axi4_lite_mosi;
   FPA_CTRL_MISO : in t_axi4_lite_miso;
   
   HEADER_CTRL_MOSI : out t_axi4_lite_mosi;
   HEADER_CTRL_MISO : in t_axi4_lite_miso;

   SFW_CTRL_MOSI : out t_axi4_lite_mosi;
   SFW_CTRL_MISO : in t_axi4_lite_miso;

   TRIGGER_CTRL_MOSI : out t_axi4_lite_mosi;
   TRIGGER_CTRL_MISO : in t_axi4_lite_miso
   
   );
end mb_model_wrapper;

architecture RTL of mb_model_wrapper is

   component mb_model
   port(
      ACLK : in STD_LOGIC;
      ARESETn : in STD_LOGIC;
      AWVALID : out STD_LOGIC_VECTOR(15 downto 0);
      AWADDR : out STD_LOGIC_VECTOR(511 downto 0);
      AWPROT : out STD_LOGIC_VECTOR(47 downto 0);
      AWREADY : in STD_LOGIC_VECTOR(15 downto 0);
      WVALID : out STD_LOGIC_VECTOR(15 downto 0);
      WREADY : in STD_LOGIC_VECTOR(15 downto 0);
      WDATA : out STD_LOGIC_VECTOR(511 downto 0);
      WSTRB : out STD_LOGIC_VECTOR(63 downto 0);
      BVALID : in STD_LOGIC_VECTOR(15 downto 0);
      BREADY : out STD_LOGIC_VECTOR(15 downto 0);
      BRESP : in STD_LOGIC_VECTOR(31 downto 0);
      ARVALID : out STD_LOGIC_VECTOR(15 downto 0);
      ARADDR : out STD_LOGIC_VECTOR(511 downto 0);
      ARPROT : out STD_LOGIC_VECTOR(47 downto 0);
      ARREADY : in STD_LOGIC_VECTOR(15 downto 0);
      RVALID : in STD_LOGIC_VECTOR(15 downto 0);
      RREADY : out STD_LOGIC_VECTOR(15 downto 0);
      RDATA : in STD_LOGIC_VECTOR(511 downto 0);
      RRESP : in STD_LOGIC_VECTOR(31 downto 0));
   end component;

--   signal ACLK_i : STD_LOGIC;
--   signal ARESETn_i : STD_LOGIC;
   signal AWVALID : STD_LOGIC_VECTOR(15 downto 0);
   signal AWADDR : STD_LOGIC_VECTOR(511 downto 0);
   signal AWPROT : STD_LOGIC_VECTOR(47 downto 0);
   signal AWREADY : STD_LOGIC_VECTOR(15 downto 0);
   signal WVALID : STD_LOGIC_VECTOR(15 downto 0);
   signal WREADY : STD_LOGIC_VECTOR(15 downto 0);
   signal WDATA : STD_LOGIC_VECTOR(511 downto 0);
   signal WSTRB : STD_LOGIC_VECTOR(63 downto 0);
   signal BVALID : STD_LOGIC_VECTOR(15 downto 0);
   signal BREADY : STD_LOGIC_VECTOR(15 downto 0);
   signal BRESP : STD_LOGIC_VECTOR(31 downto 0);
   signal ARVALID : STD_LOGIC_VECTOR(15 downto 0);
   signal ARADDR : STD_LOGIC_VECTOR(511 downto 0);
   signal ARPROT : STD_LOGIC_VECTOR(47 downto 0);
   signal ARREADY : STD_LOGIC_VECTOR(15 downto 0);
   signal RVALID : STD_LOGIC_VECTOR(15 downto 0);
   signal RREADY : STD_LOGIC_VECTOR(15 downto 0);
   signal RDATA : STD_LOGIC_VECTOR(511 downto 0);
   signal RRESP : STD_LOGIC_VECTOR(31 downto 0);
   
   

begin
   
   mb_inst : mb_model
   port map(
      ACLK => ACLK,
      ARESETn => ARESETn,
      AWVALID => AWVALID,
      AWADDR => AWADDR,
      AWPROT => AWPROT,
      AWREADY => AWREADY,
      WVALID => WVALID,
      WREADY => WREADY,
      WDATA => WDATA,
      WSTRB => WSTRB,
      BVALID => BVALID,
      BREADY => BREADY,
      BRESP => BRESP,
      ARVALID => ARVALID,
      ARADDR => ARADDR,
      ARPROT => ARPROT,
      ARREADY => ARREADY,
      RVALID => RVALID,
      RREADY => RREADY,
      RDATA => RDATA,
      RRESP => RRESP
   );
   
   --GPIO
   GPIO_MOSI.AWVALID <= AWVALID(0);
   GPIO_MOSI.AWADDR <= AWADDR(31 downto 0);
   GPIO_MOSI.AWPROT <= AWPROT(2 downto 0);
   GPIO_MOSI.WVALID <= WVALID(0);
   GPIO_MOSI.WDATA <= WDATA(31 downto 0);
   GPIO_MOSI.WSTRB <= WSTRB(3 downto 0);
   GPIO_MOSI.BREADY <= BREADY(0);
   GPIO_MOSI.ARVALID <= ARVALID(0);
   GPIO_MOSI.ARADDR <= ARADDR(31 downto 0);
   GPIO_MOSI.ARPROT <= ARPROT(2 downto 0);
   GPIO_MOSI.RREADY <= RREADY(0);
   AWREADY(0) <= GPIO_MISO.AWREADY;
   WREADY(0) <= GPIO_MISO.WREADY;
   BVALID(0) <= GPIO_MISO.BVALID;
   BRESP(1 downto 0) <= GPIO_MISO.BRESP;
   ARREADY(0) <= GPIO_MISO.ARREADY;
   RVALID(0) <= GPIO_MISO.RVALID;
   RDATA(31 downto 0) <= GPIO_MISO.RDATA;
   RRESP(1 downto 0) <= GPIO_MISO.RRESP;

   --USB_UART_MOSI
   USB_UART_MOSI.AWVALID <= AWVALID(1);
   USB_UART_MOSI.AWADDR <= AWADDR(63 downto 32);
   USB_UART_MOSI.AWPROT <= AWPROT(5 downto 3);
   USB_UART_MOSI.WVALID <= WVALID(1);
   USB_UART_MOSI.WDATA <= WDATA(63 downto 32);
   USB_UART_MOSI.WSTRB <= WSTRB(7 downto 4);
   USB_UART_MOSI.BREADY <= BREADY(1);
   USB_UART_MOSI.ARVALID <= ARVALID(1);
   USB_UART_MOSI.ARADDR <= ARADDR(63 downto 32);
   USB_UART_MOSI.ARPROT <= ARPROT(5 downto 3);
   USB_UART_MOSI.RREADY <= RREADY(1);
   AWREADY(1) <= USB_UART_MISO.AWREADY;
   WREADY(1) <= USB_UART_MISO.WREADY;
   BVALID(1) <= USB_UART_MISO.BVALID;
   BRESP(3 downto 2) <= USB_UART_MISO.BRESP;
   ARREADY(1) <= USB_UART_MISO.ARREADY;
   RVALID(1) <= USB_UART_MISO.RVALID;
   RDATA(63 downto 32) <= USB_UART_MISO.RDATA;
   RRESP(3 downto 2) <= USB_UART_MISO.RRESP;

   --CLINK_UART_MOSI
   CLINK_UART_MOSI.AWVALID <= AWVALID(2);
   CLINK_UART_MOSI.AWADDR <= AWADDR(95 downto 64);
   CLINK_UART_MOSI.AWPROT <= AWPROT(8 downto 6);
   CLINK_UART_MOSI.WVALID <= WVALID(2);
   CLINK_UART_MOSI.WDATA <= WDATA(95 downto 64);
   CLINK_UART_MOSI.WSTRB <= WSTRB(11 downto 8);
   CLINK_UART_MOSI.BREADY <= BREADY(2);
   CLINK_UART_MOSI.ARVALID <= ARVALID(2);
   CLINK_UART_MOSI.ARADDR <= ARADDR(95 downto 64);
   CLINK_UART_MOSI.ARPROT <= ARPROT(8 downto 6);
   CLINK_UART_MOSI.RREADY <= RREADY(2);
   AWREADY(2) <= CLINK_UART_MISO.AWREADY;
   WREADY(2) <= CLINK_UART_MISO.WREADY;
   BVALID(2) <= CLINK_UART_MISO.BVALID;
   BRESP(5 downto 4) <= CLINK_UART_MISO.BRESP;
   ARREADY(2) <= CLINK_UART_MISO.ARREADY;
   RVALID(2) <= CLINK_UART_MISO.RVALID;
   RDATA(95 downto 64) <= CLINK_UART_MISO.RDATA;
   RRESP(5 downto 4) <= CLINK_UART_MISO.RRESP;

   --FPGA_UART_MOSI
   FPGA_UART_MOSI.AWVALID <= AWVALID(3);
   FPGA_UART_MOSI.AWADDR <= AWADDR(127 downto 96);
   FPGA_UART_MOSI.AWPROT <= AWPROT(11 downto 9);
   FPGA_UART_MOSI.WVALID <= WVALID(3);
   FPGA_UART_MOSI.WDATA <= WDATA(127 downto 96);
   FPGA_UART_MOSI.WSTRB <= WSTRB(15 downto 12);
   FPGA_UART_MOSI.BREADY <= BREADY(3);
   FPGA_UART_MOSI.ARVALID <= ARVALID(3);
   FPGA_UART_MOSI.ARADDR <= ARADDR(127 downto 96);
   FPGA_UART_MOSI.ARPROT <= ARPROT(11 downto 9);
   FPGA_UART_MOSI.RREADY <= RREADY(3);
   AWREADY(3) <= FPGA_UART_MISO.AWREADY;
   WREADY(3) <= FPGA_UART_MISO.WREADY;
   BVALID(3) <= FPGA_UART_MISO.BVALID;
   BRESP(7 downto 6) <= FPGA_UART_MISO.BRESP;
   ARREADY(3) <= FPGA_UART_MISO.ARREADY;
   RVALID(3) <= FPGA_UART_MISO.RVALID;
   RDATA(127 downto 96) <= FPGA_UART_MISO.RDATA;
   RRESP(7 downto 6) <= FPGA_UART_MISO.RRESP;

   --OEM_UART_MOSI
   OEM_UART_MOSI.AWVALID <= AWVALID(4);
   OEM_UART_MOSI.AWADDR <= AWADDR(159 downto 128);
   OEM_UART_MOSI.AWPROT <= AWPROT(14 downto 12);
   OEM_UART_MOSI.WVALID <= WVALID(4);
   OEM_UART_MOSI.WDATA <= WDATA(159 downto 128);
   OEM_UART_MOSI.WSTRB <= WSTRB(19 downto 16);
   OEM_UART_MOSI.BREADY <= BREADY(4);
   OEM_UART_MOSI.ARVALID <= ARVALID(4);
   OEM_UART_MOSI.ARADDR <= ARADDR(159 downto 128);
   OEM_UART_MOSI.ARPROT <= ARPROT(14 downto 12);
   OEM_UART_MOSI.RREADY <= RREADY(4);
   AWREADY(4) <= OEM_UART_MISO.AWREADY;
   WREADY(4) <= OEM_UART_MISO.WREADY;
   BVALID(4) <= OEM_UART_MISO.BVALID;
   BRESP(9 downto 8) <= OEM_UART_MISO.BRESP;
   ARREADY(4) <= OEM_UART_MISO.ARREADY;
   RVALID(4) <= OEM_UART_MISO.RVALID;
   RDATA(159 downto 128) <= OEM_UART_MISO.RDATA;
   RRESP(9 downto 8) <= OEM_UART_MISO.RRESP;

   --PLEORA_UART_MOSI
   PLEORA_UART_MOSI.AWVALID <= AWVALID(5);
   PLEORA_UART_MOSI.AWADDR <= AWADDR(191 downto 160);
   PLEORA_UART_MOSI.AWPROT <= AWPROT(17 downto 15);
   PLEORA_UART_MOSI.WVALID <= WVALID(5);
   PLEORA_UART_MOSI.WDATA <= WDATA(191 downto 160);
   PLEORA_UART_MOSI.WSTRB <= WSTRB(23 downto 20);
   PLEORA_UART_MOSI.BREADY <= BREADY(5);
   PLEORA_UART_MOSI.ARVALID <= ARVALID(5);
   PLEORA_UART_MOSI.ARADDR <= ARADDR(191 downto 160);
   PLEORA_UART_MOSI.ARPROT <= ARPROT(17 downto 15);
   PLEORA_UART_MOSI.RREADY <= RREADY(5);
   AWREADY(5) <= PLEORA_UART_MISO.AWREADY;
   WREADY(5) <= PLEORA_UART_MISO.WREADY;
   BVALID(5) <= PLEORA_UART_MISO.BVALID;
   BRESP(11 downto 10) <= PLEORA_UART_MISO.BRESP;
   ARREADY(5) <= PLEORA_UART_MISO.ARREADY;
   RVALID(5) <= PLEORA_UART_MISO.RVALID;
   RDATA(191 downto 160) <= PLEORA_UART_MISO.RDATA;
   RRESP(11 downto 10) <= PLEORA_UART_MISO.RRESP;

   --XADC_MOSI
   XADC_MOSI.AWVALID <= AWVALID(6);
   XADC_MOSI.AWADDR <= AWADDR(223 downto 192);
   XADC_MOSI.AWPROT <= AWPROT(20 downto 18);
   XADC_MOSI.WVALID <= WVALID(6);
   XADC_MOSI.WDATA <= WDATA(223 downto 192);
   XADC_MOSI.WSTRB <= WSTRB(27 downto 24);
   XADC_MOSI.BREADY <= BREADY(6);
   XADC_MOSI.ARVALID <= ARVALID(6);
   XADC_MOSI.ARADDR <= ARADDR(223 downto 192);
   XADC_MOSI.ARPROT <= ARPROT(20 downto 18);
   XADC_MOSI.RREADY <= RREADY(6);
   AWREADY(6) <= XADC_MISO.AWREADY;
   WREADY(6) <= XADC_MISO.WREADY;
   BVALID(6) <= XADC_MISO.BVALID;
   BRESP(13 downto 12) <= XADC_MISO.BRESP;
   ARREADY(6) <= XADC_MISO.ARREADY;
   RVALID(6) <= XADC_MISO.RVALID;
   RDATA(223 downto 192) <= XADC_MISO.RDATA;
   RRESP(13 downto 12) <= XADC_MISO.RRESP;

   --INTC_MOSI
   INTC_MOSI.AWVALID <= AWVALID(7);
   INTC_MOSI.AWADDR <= AWADDR(255 downto 224);
   INTC_MOSI.AWPROT <= AWPROT(23 downto 21);
   INTC_MOSI.WVALID <= WVALID(7);
   INTC_MOSI.WDATA <= WDATA(255 downto 224);
   INTC_MOSI.WSTRB <= WSTRB(31 downto 28);
   INTC_MOSI.BREADY <= BREADY(7);
   INTC_MOSI.ARVALID <= ARVALID(7);
   INTC_MOSI.ARADDR <= ARADDR(255 downto 224);
   INTC_MOSI.ARPROT <= ARPROT(23 downto 21);
   INTC_MOSI.RREADY <= RREADY(7);
   AWREADY(7) <= INTC_MISO.AWREADY;
   WREADY(7) <= INTC_MISO.WREADY;
   BVALID(7) <= INTC_MISO.BVALID;
   BRESP(15 downto 14) <= INTC_MISO.BRESP;
   ARREADY(7) <= INTC_MISO.ARREADY;
   RVALID(7) <= INTC_MISO.RVALID;
   RDATA(255 downto 224) <= INTC_MISO.RDATA;
   RRESP(15 downto 14) <= INTC_MISO.RRESP;

   --AEC_CTRL_MOSI
   AEC_CTRL_MOSI.AWVALID <= AWVALID(8);
   AEC_CTRL_MOSI.AWADDR <= AWADDR(287 downto 256);
   AEC_CTRL_MOSI.AWPROT <= AWPROT(26 downto 24);
   AEC_CTRL_MOSI.WVALID <= WVALID(8);
   AEC_CTRL_MOSI.WDATA <= WDATA(287 downto 256);
   AEC_CTRL_MOSI.WSTRB <= WSTRB(35 downto 32);
   AEC_CTRL_MOSI.BREADY <= BREADY(8);
   AEC_CTRL_MOSI.ARVALID <= ARVALID(8);
   AEC_CTRL_MOSI.ARADDR <= ARADDR(287 downto 256);
   AEC_CTRL_MOSI.ARPROT <= ARPROT(26 downto 24);
   AEC_CTRL_MOSI.RREADY <= RREADY(8);
   AWREADY(8) <= AEC_CTRL_MISO.AWREADY;
   WREADY(8) <= AEC_CTRL_MISO.WREADY;
   BVALID(8) <= AEC_CTRL_MISO.BVALID;
   BRESP(17 downto 16) <= AEC_CTRL_MISO.BRESP;
   ARREADY(8) <= AEC_CTRL_MISO.ARREADY;
   RVALID(8) <= AEC_CTRL_MISO.RVALID;
   RDATA(287 downto 256) <= AEC_CTRL_MISO.RDATA;
   RRESP(17 downto 16) <= AEC_CTRL_MISO.RRESP;

   --BPR_CTRL_MOSI
   BPR_CTRL_MOSI.AWVALID <= AWVALID(9);
   BPR_CTRL_MOSI.AWADDR <= AWADDR(319 downto 288);
   BPR_CTRL_MOSI.AWPROT <= AWPROT(29 downto 27);
   BPR_CTRL_MOSI.WVALID <= WVALID(9);
   BPR_CTRL_MOSI.WDATA <= WDATA(319 downto 288);
   BPR_CTRL_MOSI.WSTRB <= WSTRB(39 downto 36);
   BPR_CTRL_MOSI.BREADY <= BREADY(9);
   BPR_CTRL_MOSI.ARVALID <= ARVALID(9);
   BPR_CTRL_MOSI.ARADDR <= ARADDR(319 downto 288);
   BPR_CTRL_MOSI.ARPROT <= ARPROT(29 downto 27);
   BPR_CTRL_MOSI.RREADY <= RREADY(9);
   AWREADY(9) <= BPR_CTRL_MISO.AWREADY;
   WREADY(9) <= BPR_CTRL_MISO.WREADY;
   BVALID(9) <= BPR_CTRL_MISO.BVALID;
   BRESP(19 downto 18) <= BPR_CTRL_MISO.BRESP;
   ARREADY(9) <= BPR_CTRL_MISO.ARREADY;
   RVALID(9) <= BPR_CTRL_MISO.RVALID;
   RDATA(319 downto 288) <= BPR_CTRL_MISO.RDATA;
   RRESP(19 downto 18) <= BPR_CTRL_MISO.RRESP;

   --CAL_CTRL_MOSI
   CAL_CTRL_MOSI.AWVALID <= AWVALID(10);
   CAL_CTRL_MOSI.AWADDR <= AWADDR(351 downto 320);
   CAL_CTRL_MOSI.AWPROT <= AWPROT(32 downto 30);
   CAL_CTRL_MOSI.WVALID <= WVALID(10);
   CAL_CTRL_MOSI.WDATA <= WDATA(351 downto 320);
   CAL_CTRL_MOSI.WSTRB <= WSTRB(43 downto 40);
   CAL_CTRL_MOSI.BREADY <= BREADY(10);
   CAL_CTRL_MOSI.ARVALID <= ARVALID(10);
   CAL_CTRL_MOSI.ARADDR <= ARADDR(351 downto 320);
   CAL_CTRL_MOSI.ARPROT <= ARPROT(32 downto 30);
   CAL_CTRL_MOSI.RREADY <= RREADY(10);
   AWREADY(10) <= CAL_CTRL_MISO.AWREADY;
   WREADY(10) <= CAL_CTRL_MISO.WREADY;
   BVALID(10) <= CAL_CTRL_MISO.BVALID;
   BRESP(21 downto 20) <= CAL_CTRL_MISO.BRESP;
   ARREADY(10) <= CAL_CTRL_MISO.ARREADY;
   RVALID(10) <= CAL_CTRL_MISO.RVALID;
   RDATA(351 downto 320) <= CAL_CTRL_MISO.RDATA;
   RRESP(21 downto 20) <= CAL_CTRL_MISO.RRESP;

   --EXPTIME_CTRL_MOSI
   EXPTIME_CTRL_MOSI.AWVALID <= AWVALID(11);
   EXPTIME_CTRL_MOSI.AWADDR <= AWADDR(383 downto 352);
   EXPTIME_CTRL_MOSI.AWPROT <= AWPROT(35 downto 33);
   EXPTIME_CTRL_MOSI.WVALID <= WVALID(11);
   EXPTIME_CTRL_MOSI.WDATA <= WDATA(383 downto 352);
   EXPTIME_CTRL_MOSI.WSTRB <= WSTRB(47 downto 44);
   EXPTIME_CTRL_MOSI.BREADY <= BREADY(11);
   EXPTIME_CTRL_MOSI.ARVALID <= ARVALID(11);
   EXPTIME_CTRL_MOSI.ARADDR <= ARADDR(383 downto 352);
   EXPTIME_CTRL_MOSI.ARPROT <= ARPROT(35 downto 33);
   EXPTIME_CTRL_MOSI.RREADY <= RREADY(11);
   AWREADY(11) <= EXPTIME_CTRL_MISO.AWREADY;
   WREADY(11) <= EXPTIME_CTRL_MISO.WREADY;
   BVALID(11) <= EXPTIME_CTRL_MISO.BVALID;
   BRESP(23 downto 22) <= EXPTIME_CTRL_MISO.BRESP;
   ARREADY(11) <= EXPTIME_CTRL_MISO.ARREADY;
   RVALID(11) <= EXPTIME_CTRL_MISO.RVALID;
   RDATA(383 downto 352) <= EXPTIME_CTRL_MISO.RDATA;
   RRESP(23 downto 22) <= EXPTIME_CTRL_MISO.RRESP;

   --FPA_CTRL_MOSI
   FPA_CTRL_MOSI.AWVALID <= AWVALID(12);
   FPA_CTRL_MOSI.AWADDR <= AWADDR(415 downto 384);
   FPA_CTRL_MOSI.AWPROT <= AWPROT(38 downto 36);
   FPA_CTRL_MOSI.WVALID <= WVALID(12);
   FPA_CTRL_MOSI.WDATA <= WDATA(415 downto 384);
   FPA_CTRL_MOSI.WSTRB <= WSTRB(51 downto 48);
   FPA_CTRL_MOSI.BREADY <= BREADY(12);
   FPA_CTRL_MOSI.ARVALID <= ARVALID(12);
   FPA_CTRL_MOSI.ARADDR <= ARADDR(415 downto 384);
   FPA_CTRL_MOSI.ARPROT <= ARPROT(38 downto 36);
   FPA_CTRL_MOSI.RREADY <= RREADY(12);
   AWREADY(12) <= FPA_CTRL_MISO.AWREADY;
   WREADY(12) <= FPA_CTRL_MISO.WREADY;
   BVALID(12) <= FPA_CTRL_MISO.BVALID;
   BRESP(25 downto 24) <= FPA_CTRL_MISO.BRESP;
   ARREADY(12) <= FPA_CTRL_MISO.ARREADY;
   RVALID(12) <= FPA_CTRL_MISO.RVALID;
   RDATA(415 downto 384) <= FPA_CTRL_MISO.RDATA;
   RRESP(25 downto 24) <= FPA_CTRL_MISO.RRESP;

   --HEADER_CTRL_MOSI
   HEADER_CTRL_MOSI.AWVALID <= AWVALID(13);
   HEADER_CTRL_MOSI.AWADDR <= AWADDR(447 downto 416);
   HEADER_CTRL_MOSI.AWPROT <= AWPROT(41 downto 39);
   HEADER_CTRL_MOSI.WVALID <= WVALID(13);
   HEADER_CTRL_MOSI.WDATA <= WDATA(447 downto 416);
   HEADER_CTRL_MOSI.WSTRB <= WSTRB(55 downto 52);
   HEADER_CTRL_MOSI.BREADY <= BREADY(13);
   HEADER_CTRL_MOSI.ARVALID <= ARVALID(13);
   HEADER_CTRL_MOSI.ARADDR <= ARADDR(447 downto 416);
   HEADER_CTRL_MOSI.ARPROT <= ARPROT(41 downto 39);
   HEADER_CTRL_MOSI.RREADY <= RREADY(13);
   AWREADY(13) <= HEADER_CTRL_MISO.AWREADY;
   WREADY(13) <= HEADER_CTRL_MISO.WREADY;
   BVALID(13) <= HEADER_CTRL_MISO.BVALID;
   BRESP(27 downto 26) <= HEADER_CTRL_MISO.BRESP;
   ARREADY(13) <= HEADER_CTRL_MISO.ARREADY;
   RVALID(13) <= HEADER_CTRL_MISO.RVALID;
   RDATA(447 downto 416) <= HEADER_CTRL_MISO.RDATA;
   RRESP(27 downto 26) <= HEADER_CTRL_MISO.RRESP;

   --SFW_CTRL_MOSI
   SFW_CTRL_MOSI.AWVALID <= AWVALID(14);
   SFW_CTRL_MOSI.AWADDR <= AWADDR(479 downto 448);
   SFW_CTRL_MOSI.AWPROT <= AWPROT(44 downto 42);
   SFW_CTRL_MOSI.WVALID <= WVALID(14);
   SFW_CTRL_MOSI.WDATA <= WDATA(479 downto 448);
   SFW_CTRL_MOSI.WSTRB <= WSTRB(59 downto 56);
   SFW_CTRL_MOSI.BREADY <= BREADY(14);
   SFW_CTRL_MOSI.ARVALID <= ARVALID(14);
   SFW_CTRL_MOSI.ARADDR <= ARADDR(479 downto 448);
   SFW_CTRL_MOSI.ARPROT <= ARPROT(44 downto 42);
   SFW_CTRL_MOSI.RREADY <= RREADY(14);
   AWREADY(14) <= SFW_CTRL_MISO.AWREADY;
   WREADY(14) <= SFW_CTRL_MISO.WREADY;
   BVALID(14) <= SFW_CTRL_MISO.BVALID;
   BRESP(29 downto 28) <= SFW_CTRL_MISO.BRESP;
   ARREADY(14) <= SFW_CTRL_MISO.ARREADY;
   RVALID(14) <= SFW_CTRL_MISO.RVALID;
   RDATA(479 downto 448) <= SFW_CTRL_MISO.RDATA;
   RRESP(29 downto 28) <= SFW_CTRL_MISO.RRESP;

   --SFW_CTRL_MOSI
   TRIGGER_CTRL_MOSI.AWVALID <= AWVALID(15);
   TRIGGER_CTRL_MOSI.AWADDR <= AWADDR(511 downto 480);
   TRIGGER_CTRL_MOSI.AWPROT <= AWPROT(47 downto 45);
   TRIGGER_CTRL_MOSI.WVALID <= WVALID(15);
   TRIGGER_CTRL_MOSI.WDATA <= WDATA(511 downto 480);
   TRIGGER_CTRL_MOSI.WSTRB <= WSTRB(63 downto 60);
   TRIGGER_CTRL_MOSI.BREADY <= BREADY(15);
   TRIGGER_CTRL_MOSI.ARVALID <= ARVALID(15);
   TRIGGER_CTRL_MOSI.ARADDR <= ARADDR(511 downto 480);
   TRIGGER_CTRL_MOSI.ARPROT <= ARPROT(47 downto 45);
   TRIGGER_CTRL_MOSI.RREADY <= RREADY(15);
   AWREADY(15) <= TRIGGER_CTRL_MISO.AWREADY;
   WREADY(15) <= TRIGGER_CTRL_MISO.WREADY;
   BVALID(15) <= TRIGGER_CTRL_MISO.BVALID;
   BRESP(31 downto 30) <= TRIGGER_CTRL_MISO.BRESP;
   ARREADY(15) <= TRIGGER_CTRL_MISO.ARREADY;
   RVALID(15) <= TRIGGER_CTRL_MISO.RVALID;
   RDATA(511 downto 480) <= TRIGGER_CTRL_MISO.RDATA;
   RRESP(31 downto 30) <= TRIGGER_CTRL_MISO.RRESP;

end RTL;