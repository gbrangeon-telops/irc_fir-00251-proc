--******************************************************************************
-- Destination: 
--
--	File: Proxy_define.vhd
-- Hierarchy: Package file
-- Use: 
--	Project: IRCDEV
--	By: Edem Nofodjie
-- Date: 22 october 2009	  
--
--******************************************************************************
--Description
--******************************************************************************
-- 1- Defines the global variables 
-- 2- Defines the project function
--******************************************************************************


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use work.fpa_common_pkg.all;
use work.fpa_define.all;  

package Proxy_define is
   
   --------------------------------------------
   -- PROJET: definition
   --------------------------------------------   
   constant DEFINE_PROXY                 : std_logic_vector(2 downto 0) := PROXY_BB1920D;
   constant PROG_FREE_RUNNING_TRIG       : std_logic := '0';   -- � '1', cette constante dit que les trigs n'ont pas besoin d'�tre arr�t� lorsqu'on programme le d�tecteur
   constant FPA_INTF_CLK_RATE_MHZ        : integer := 100;     --  FPA_INTF_CLK_RATE en MHz
   constant BB1920D_INT_TIME_MIN_US          : integer := 1; 
   constant BB1920D_MASTER_CLK_RATE_MHZ      : integer := 80;      --
   constant FPA_XTRA_IMAGE_NUM_TO_SKIP   : integer := 1; -- pour le pelicanD, chaque appel de FPA_SendConfigGC() d�clenche l'envoi d'une config op�rationnelle au proxy qui sera pr�c�d� et suivi d'au moins FPA_XTRA_IMAGE_NUM_TO_SKIP prog trig.  
   --constant PROXY_CLINK_CHANNEL_NUM      : integer := DEFINE_FPA_CLINK_CHANNEL_NUM;     -- Number of channels in the Camera Link interface with the proxy 
   --constant PROXY_CLINK_CLK_1X_PERIOD_NS : real    := 12.5;  -- CLINK IN est � 80MHz ns pour les BB1920D
   --------------------------------------------
   --  modes diag
   --------------------------------------------
   -- D comme diag mais en fait pour laisser les valeurs inf�rieurs au
   constant TELOPS_DIAG_CNST             : std_logic_vector(7 downto 0):= x"D1";  -- mode diag constant
   constant TELOPS_DIAG_DEGR             : std_logic_vector(7 downto 0):= x"D2";  -- mode diag degrad� pour la prod
   constant TELOPS_DIAG_DEGR_DYN         : std_logic_vector(7 downto 0):= x"D3";  -- mode diag degrad� dynamique pour FAU
   
   --------------------------------------------
   -- FPA : Nombre d'ADCs sur le FPA
   -------------------------------------------- 
   constant NUMBER_TAPS                  : natural := 1;
   
   ----------------------------------------------
   -- FPA 
   ---------------------------------------------- 
   constant BB1920D_GAIN_0                   : std_logic_vector(7 downto 0) := x"00";
   constant BB1920D_GAIN_1                   : std_logic_vector(7 downto 0) := x"02";
   constant BB1920D_ITR                      : std_logic_vector(7 downto 0) := x"00";
   constant BB1920D_IWR                      : std_logic_vector(7 downto 0) := x"01";
   constant BB1920D_PIX_RES_15B              : std_logic_vector(1 downto 0) := "00";
   constant BB1920D_PIX_RES_14B              : std_logic_vector(1 downto 0) := "01";
   constant BB1920D_PIX_RES_13B              : std_logic_vector(1 downto 0) := "10";
   constant FPA_INT_FBK_AVAILABLE        : std_logic := '1';
   constant BB1920D_FSYNC_HIGH_TIME_US       : integer := 5;     -- duree de FSYNC en usec
   constant BB1920D_POWER_WAIT_US            : integer := 2_000_000;  -- duree d'attente apr�s allumage en usec. selon la doc, le proxy prend 1 sec. Pour plus de securit�, j'en mets 2
   constant BB1920D_TEMP_TRIG_PERIOD_US      : integer := 1_000_000;  -- le trig de lecture de la temperature a une periode de 1sec pour ne pas submerger le proxy
   
   -- commandes
   constant BB1920D_CMD_OVERHEAD_BYTES_NUM   : integer := 6; -- nombre de bytes de l'overhead (header, CommandID, length, Checksum)
   constant BB1920D_LONGEST_CMD_BYTES_NUM    : integer := 32; -- longueur maximale en byte de la config d'un bb1920D (incluant le header, checksum etc). Ce nombre doit �tre inf�rieur � 64 � cause d'un fifo dans le copieur
   constant BB1920D_SERIAL_BAUD_RATE         : integer := 921_600; -- baud rate utilis� pour Scd (utilis� juste pour generateur de delai)
   constant BB1920D_COM_RESP_HDER            : std_logic_vector(7 downto 0)  := x"55";
   constant BB1920D_COM_RESP_FAILURE_ID      : std_logic_vector(15 downto 0) := x"FFFF";
   constant BB1920D_CMD_HDER                 : std_logic_vector(7 downto 0)  := x"AA";
   
   -- serial int time cmd
   constant BB1920D_INT_CMD_ID               : std_logic_vector(15 downto 0) := x"8001";
   constant BB1920D_INT_CMD_DLEN             : std_logic_vector(15 downto 0) := x"0006";
   
   -- serial operational cmd
   constant BB1920D_OP_CMD_ID                : std_logic_vector(15 downto 0) := x"8002";
   
   -- serial diag cmd                                                        
   constant BB1920D_DIAG_CMD_ID              : std_logic_vector(15 downto 0) := x"8004";
   
   -- serial temperature read cmd
   constant BB1920D_TEMP_CMD_ID              : std_logic_vector(15 downto 0) := x"8021";
   
   -- partition de la ram de cfg serielle (la partie d'ecriture reserv�e � la config serielle a une plage d'adresse < 255)
   constant BB1920D_OP_CMD_RAM_BASE_ADD      : integer  := 0;    -- adresse de base o� est log�e la commande operationnelle en ram
   constant BB1920D_INT_CMD_RAM_BASE_ADD     : integer  := 64;   -- adresse de base o� est log�e la commande du temps d'integration en ram
   constant BB1920D_DIAG_CMD_RAM_BASE_ADD    : integer  := 128;
   constant BB1920D_TEMP_CMD_RAM_BASE_ADD    : integer  := 192;
   
   -- adresse de base de la zone securis�e
   constant BB1920D_CMD_SECUR_RAM_BASE_ADD   : integer  := 1024; -- adresse o� se retrouve la commande copi�e dans la zone securisee
   
   -- quelques constantes 
   constant SERIAL_CFG_END_ADD           : std_logic_vector(7 downto 0) := x"FC"; -- adresse de fin d'envoi de la config serielle
   constant SERIAL_CFG_COPIER_START_DLY  : integer := 10; -- delai ajust� par simulation pour eviter corruption de config dans la RAM
   constant SERIAL_CFG_COPIER_END_DLY    : integer := 10; -- delai ajust� par simulation pour eviter corruption de config dans la RAM
   
   ----------------------------------------------
   -- Calculs 
   ---------------------------------------------- 
   constant BB1920D_FSYNC_HIGH_TIME_FACTOR     : integer := integer(FPA_INTF_CLK_RATE_MHZ*BB1920D_FSYNC_HIGH_TIME_US);
   constant BB1920D_POWER_WAIT_FACTOR          : integer := integer(FPA_INTF_CLK_RATE_MHZ*BB1920D_POWER_WAIT_US);
   constant BB1920D_SERIAL_TX_CLK_FACTOR       : integer := integer((FPA_INTF_CLK_RATE_MHZ*1E6)/BB1920D_SERIAL_BAUD_RATE); -- utilis� juste pour generateur de delai
   constant BB1920D_OP_INT_TIME_DEFAULT_FACTOR : integer := integer(real(BB1920D_MASTER_CLK_RATE_MHZ)*(0.5*real(BB1920D_INT_TIME_MIN_US))); --
   constant BB1920D_TEMP_TRIG_PERIOD_FACTOR    : integer := integer(FPA_INTF_CLK_RATE_MHZ*BB1920D_TEMP_TRIG_PERIOD_US);
   
   constant BB1920D_EXP_TIME_CONV_DENOMINATOR_BIT_POS : natural := 26;  -- log2 de BB1920D_EXP_TIME_CONV_DENOMINATOR  
   constant BB1920D_EXP_TIME_CONV_DENOMINATOR  : integer := 2**BB1920D_EXP_TIME_CONV_DENOMINATOR_BIT_POS;
   constant BB1920D_EXP_TIME_CONV_NUMERATOR    : unsigned(BB1920D_EXP_TIME_CONV_DENOMINATOR_BIT_POS-1 downto 0):= to_unsigned((4*(2**BB1920D_EXP_TIME_CONV_DENOMINATOR_BIT_POS))/5, BB1920D_EXP_TIME_CONV_DENOMINATOR_BIT_POS);     -- (80 x 2^26 )/100
   constant DEFINE_DIAG_DATA_CLK_FACTOR    : integer := integer(ceil(real(FPA_INTF_CLK_RATE_MHZ * 1000) / real(DEFINE_DIAG_CLK_RATE_MAX_KHZ)));  
   
   
   
   ---------------------------------------------------------------------------------								
   -- Configuration regroupant les �l�ments vraiment propres au d�tecteur
   ---------------------------------------------------------------------------------
   -- bb1920D integration
   type bb1920D_int_cfg_type is
   record
      bb1920D_int_time            : unsigned(23 downto 0);  --! temps d'integration en coups de 80Mhz
      diag_int_time           : unsigned(24 downto 0);  --! temps d'integration en coups de 100Mhz
      bb1920D_int_indx            : std_logic_vector(7 downto 0);
   end record;
   
   -- bb1920D operationnelle
   type bb1920D_op_cfg_type is
   record  
      bb1920D_xstart              : unsigned(10 downto 0); 
      bb1920D_ystart              : unsigned(10 downto 0);
      bb1920D_xsize               : unsigned(10 downto 0);
      bb1920D_ysize               : unsigned(10 downto 0);
      bb1920D_gain                : std_logic_vector(7 downto 0);
      bb1920D_out_chn             : std_logic;
      bb1920D_diode_bias          : std_logic_vector(3 downto 0);
      bb1920D_int_mode            : std_logic_vector(7 downto 0);
      bb1920D_boost_mode          : std_logic;
      bb1920D_pix_res             : std_logic_vector(1 downto 0);
      bb1920D_frame_period_min    : unsigned(23 downto 0); 
      cfg_num                 : unsigned(7 downto 0);      
   end record;
   
   -- bb1920D video synthetic
   type bb1920D_diag_cfg_type is
   record
      bb1920D_bit_pattern         : std_logic_vector(2 downto 0);   
   end record;
   
   -- bb1920D temperature
   type bb1920D_temp_cfg_type is
   record
      bb1920D_temp_read_num       : unsigned(7 downto 0);
   end record; 
   
   -- bb1920D misc                 --  quelques valeurs propres au PelicanD (-- se reporter aux figures 1 et 2 et 4 des pages 13, 15 et 19 du doument Communication protocol appendix A5 (SPEC. NO: DPS3008) dans le dossier du pelicanD)                                
   type bb1920D_misc_cfg_type is
   record
      bb1920D_fig1_or_fig2_t6_dly : unsigned(15 downto 0);
      bb1920D_fig4_t1_dly         : unsigned(15 downto 0);
      bb1920D_fig4_t2_dly         : unsigned(15 downto 0);
      bb1920D_fig4_t6_dly         : unsigned(15 downto 0);
      bb1920D_fig4_t3_dly         : unsigned(15 downto 0);
      bb1920D_fig4_t5_dly         : unsigned(15 downto 0);
      bb1920D_fig4_t4_dly         : unsigned(15 downto 0);
      bb1920D_fig1_or_fig2_t5_dly : unsigned(15 downto 0);
      bb1920D_fig1_or_fig2_t4_dly : unsigned(15 downto 0);
      bb1920D_xsize_div2          : unsigned(9 downto 0);
   end record;
   
   ------------------------------------------------								
   -- Configuration du Bloc FPA_interface
   ------------------------------------------------
   type fpa_intf_cfg_type is
   record     
      cmd_to_update_id     : std_logic_vector(15 downto 0); -- cet ide permet de saoir quelle partie de la commande rentrante est � mettre � jour. Important pour regler bugs
      comn                 : fpa_comn_cfg_type;   -- partie commune (utilis�e par les modules communs)
      bb1920D_op               : bb1920D_op_cfg_type;     -- tout changement dans bb1920D_op entraine la programmation du detecteur (commnde operationnelle)
      bb1920D_int              : bb1920D_int_cfg_type;    -- tout changement dans bb1920D_int entraine la programmation du detecteur (commnde temps d'int�gration)
      bb1920D_diag             : bb1920D_diag_cfg_type;   -- tout changement dans bb1920D_diag entraine la programmation du detecteur (commnde PE Syntehtique)
      bb1920D_temp             : bb1920D_temp_cfg_type;   -- tout changement dans bb1920D_temp entraine la programmation du detecteur (commnde temperature read)  
      bb1920D_misc             : bb1920D_misc_cfg_type;   -- les changements dans bb1920D_misc ne font pas programmer le detecteur
      fpa_serdes_lval_num  : unsigned(10 downto 0);   -- pour la calibration des serdes d'entr�e
      fpa_serdes_lval_len  : unsigned(10 downto 0);   -- pour la calibration des serdes d'entr�e
      int_time             : unsigned(31 downto 0);   -- temps d'integration actuellement utilis� en coups de MCLK. Sert juste � generer un statut.
   end record;    
   
   ----------------------------------------------								
   -- Type hder_param
   ----------------------------------------------
   type hder_param_type is
   record
      exp_time            : unsigned(31 downto 0); -- temps d'integration en coups de 100 MHz
      frame_id            : unsigned(31 downto 0);
      sensor_temp_raw     : std_logic_vector(15 downto 0);
      exp_index           : unsigned(7 downto 0);
      rdy                 : std_logic;                     -- pulse signifiant que les parametres du header sont pr�ts
   end record;
   
   
   ----------------------------------------------								
   -- Type diag_data_ofs_type
   ----------------------------------------------
   --type diag_data_ofs_type is array (1 to 9) of natural range 0 to ((2**16)*9)/XSIZE_MAX; -- (1 to 9) pour accommoder 4 ou 8 taps
   
   
   ----------------------------------------------
   -- quues fontions                                    
   ----------------------------------------------
   --function to_diag_data_ofs return diag_data_ofs_type;
   --function to_fpa_word_func(a:fpa_intf_cfg_type) return fpa_word_type;

end Proxy_define;

package body Proxy_define is
   
   ---
   -- function to_diag_data_ofs return diag_data_ofs_type is
      -- variable y  : diag_data_ofs_type;
      -- variable ii : integer range 1 to 9;
      
   -- begin
      -- for ii in 1 to 9 loop    
         -- y(ii) := (ii - 1)*DIAG_DATA_INC;
      -- end loop;   
      -- return y;                 
   -- end to_diag_data_ofs; 
   
end package body Proxy_define; 
